module MIPS_tb();

endmodule