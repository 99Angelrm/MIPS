module MIPS ();

endmodule